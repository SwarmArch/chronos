ARG_WIDTH 16

core des_core 7
core des_enqueuer 1
