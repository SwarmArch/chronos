ARG_WIDTH 1

core sssp_hls 8
