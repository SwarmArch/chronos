
parameter APP_NAME = "color";
parameter RISCV = 0;

parameter ARG_WIDTH = 80;

parameter RW_WIDTH = 256;
parameter DATA_WIDTH = 32;

parameter LOG_N_SUB_TYPES = 1;


`define RO_WORKER color_worker
`define RW_WORKER color_rw
