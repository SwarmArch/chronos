# ARG_WIDTH has to be a multiple of 32
ARG_WIDTH 128
 
APP_ID 256
RISCV_APP sssp

mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
