ARG_WIDTH 64
RISCV_APP maxflow

mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
