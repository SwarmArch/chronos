ARG_WIDTH 64
RISCV_APP sssp

mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
mt_core riscv_core 1
