ARG_WIDTH 16
APP_ID 1

core des_core 7
core des_enqueuer 1
