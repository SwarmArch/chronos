ARG_WIDTH 64

core visit_vertex 8 
core terminate_core 1 
mt_core queue_vertex 16
