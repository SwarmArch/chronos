ARG_WIDTH 32
# core module_name num_cores 
core color 8 all_tasks
