ARG_WIDTH 1
APP_ID 0

core sssp_core 8
