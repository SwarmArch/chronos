ARG_WIDTH 32
APP_ID 4
# core module_name num_cores 
core color 8 all_tasks
