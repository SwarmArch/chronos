ARG_WIDTH 1

core sssp_core 8
