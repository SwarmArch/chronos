ARG_WIDTH 64
DATA_WIDTH 64
APP_ID 3

# core module_name num_cores 
core maxflow 8 all_tasks
