ARG_WIDTH 64
# core module_name num_cores 
core maxflow 8 all_tasks
